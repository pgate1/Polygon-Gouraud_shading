
/*Produced by sfl2vl, IP ARCH, Inc. Sun Jul 14 18:45:30 2019
 Licensed to :EVALUATION USER*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module inv_table ( p_reset , m_clock , dout , read , adrs );
  input p_reset, m_clock;
  wire p_reset, m_clock;
  output [15:0] dout;
  wire [15:0] dout;
  input read;
  wire read;
  input [9:0] adrs;
  wire [9:0] adrs;
  reg [15:0] dout_reg;
  reg [15:0] cells [0:1023];

   assign  dout = dout_reg;
always @(posedge m_clock or posedge p_reset)
  begin
if (p_reset)
     dout_reg <= 16'b0000000000000000;
else if ((read)) 
      dout_reg <= (cells[adrs]);
end
initial begin
    cells[0] = 16'b0000000000000000;
    cells[1] = 16'b0111111111111111;
    cells[2] = 16'b0100000000000000;
    cells[3] = 16'b0010101010101010;
    cells[4] = 16'b0010000000000000;
    cells[5] = 16'b0001100110011001;
    cells[6] = 16'b0001010101010101;
    cells[7] = 16'b0001001001001001;
    cells[8] = 16'b0001000000000000;
    cells[9] = 16'b0000111000111000;
    cells[10] = 16'b0000110011001100;
    cells[11] = 16'b0000101110100010;
    cells[12] = 16'b0000101010101010;
    cells[13] = 16'b0000100111011000;
    cells[14] = 16'b0000100100100100;
    cells[15] = 16'b0000100010001000;
    cells[16] = 16'b0000100000000000;
    cells[17] = 16'b0000011110000111;
    cells[18] = 16'b0000011100011100;
    cells[19] = 16'b0000011010111100;
    cells[20] = 16'b0000011001100110;
    cells[21] = 16'b0000011000011000;
    cells[22] = 16'b0000010111010001;
    cells[23] = 16'b0000010110010000;
    cells[24] = 16'b0000010101010101;
    cells[25] = 16'b0000010100011110;
    cells[26] = 16'b0000010011101100;
    cells[27] = 16'b0000010010111101;
    cells[28] = 16'b0000010010010010;
    cells[29] = 16'b0000010001101001;
    cells[30] = 16'b0000010001000100;
    cells[31] = 16'b0000010000100001;
    cells[32] = 16'b0000010000000000;
    cells[33] = 16'b0000001111100000;
    cells[34] = 16'b0000001111000011;
    cells[35] = 16'b0000001110101000;
    cells[36] = 16'b0000001110001110;
    cells[37] = 16'b0000001101110101;
    cells[38] = 16'b0000001101011110;
    cells[39] = 16'b0000001101001000;
    cells[40] = 16'b0000001100110011;
    cells[41] = 16'b0000001100011111;
    cells[42] = 16'b0000001100001100;
    cells[43] = 16'b0000001011111010;
    cells[44] = 16'b0000001011101000;
    cells[45] = 16'b0000001011011000;
    cells[46] = 16'b0000001011001000;
    cells[47] = 16'b0000001010111001;
    cells[48] = 16'b0000001010101010;
    cells[49] = 16'b0000001010011100;
    cells[50] = 16'b0000001010001111;
    cells[51] = 16'b0000001010000010;
    cells[52] = 16'b0000001001110110;
    cells[53] = 16'b0000001001101010;
    cells[54] = 16'b0000001001011110;
    cells[55] = 16'b0000001001010011;
    cells[56] = 16'b0000001001001001;
    cells[57] = 16'b0000001000111110;
    cells[58] = 16'b0000001000110100;
    cells[59] = 16'b0000001000101011;
    cells[60] = 16'b0000001000100010;
    cells[61] = 16'b0000001000011001;
    cells[62] = 16'b0000001000010000;
    cells[63] = 16'b0000001000001000;
    cells[64] = 16'b0000001000000000;
    cells[65] = 16'b0000000111111000;
    cells[66] = 16'b0000000111110000;
    cells[67] = 16'b0000000111101001;
    cells[68] = 16'b0000000111100001;
    cells[69] = 16'b0000000111011010;
    cells[70] = 16'b0000000111010100;
    cells[71] = 16'b0000000111001101;
    cells[72] = 16'b0000000111000111;
    cells[73] = 16'b0000000111000000;
    cells[74] = 16'b0000000110111010;
    cells[75] = 16'b0000000110110100;
    cells[76] = 16'b0000000110101111;
    cells[77] = 16'b0000000110101001;
    cells[78] = 16'b0000000110100100;
    cells[79] = 16'b0000000110011110;
    cells[80] = 16'b0000000110011001;
    cells[81] = 16'b0000000110010100;
    cells[82] = 16'b0000000110001111;
    cells[83] = 16'b0000000110001010;
    cells[84] = 16'b0000000110000110;
    cells[85] = 16'b0000000110000001;
    cells[86] = 16'b0000000101111101;
    cells[87] = 16'b0000000101111000;
    cells[88] = 16'b0000000101110100;
    cells[89] = 16'b0000000101110000;
    cells[90] = 16'b0000000101101100;
    cells[91] = 16'b0000000101101000;
    cells[92] = 16'b0000000101100100;
    cells[93] = 16'b0000000101100000;
    cells[94] = 16'b0000000101011100;
    cells[95] = 16'b0000000101011000;
    cells[96] = 16'b0000000101010101;
    cells[97] = 16'b0000000101010001;
    cells[98] = 16'b0000000101001110;
    cells[99] = 16'b0000000101001010;
    cells[100] = 16'b0000000101000111;
    cells[101] = 16'b0000000101000100;
    cells[102] = 16'b0000000101000001;
    cells[103] = 16'b0000000100111110;
    cells[104] = 16'b0000000100111011;
    cells[105] = 16'b0000000100111000;
    cells[106] = 16'b0000000100110101;
    cells[107] = 16'b0000000100110010;
    cells[108] = 16'b0000000100101111;
    cells[109] = 16'b0000000100101100;
    cells[110] = 16'b0000000100101001;
    cells[111] = 16'b0000000100100111;
    cells[112] = 16'b0000000100100100;
    cells[113] = 16'b0000000100100001;
    cells[114] = 16'b0000000100011111;
    cells[115] = 16'b0000000100011100;
    cells[116] = 16'b0000000100011010;
    cells[117] = 16'b0000000100011000;
    cells[118] = 16'b0000000100010101;
    cells[119] = 16'b0000000100010011;
    cells[120] = 16'b0000000100010001;
    cells[121] = 16'b0000000100001110;
    cells[122] = 16'b0000000100001100;
    cells[123] = 16'b0000000100001010;
    cells[124] = 16'b0000000100001000;
    cells[125] = 16'b0000000100000110;
    cells[126] = 16'b0000000100000100;
    cells[127] = 16'b0000000100000010;
    cells[128] = 16'b0000000100000000;
    cells[129] = 16'b0000000011111110;
    cells[130] = 16'b0000000011111100;
    cells[131] = 16'b0000000011111010;
    cells[132] = 16'b0000000011111000;
    cells[133] = 16'b0000000011110110;
    cells[134] = 16'b0000000011110100;
    cells[135] = 16'b0000000011110010;
    cells[136] = 16'b0000000011110000;
    cells[137] = 16'b0000000011101111;
    cells[138] = 16'b0000000011101101;
    cells[139] = 16'b0000000011101011;
    cells[140] = 16'b0000000011101010;
    cells[141] = 16'b0000000011101000;
    cells[142] = 16'b0000000011100110;
    cells[143] = 16'b0000000011100101;
    cells[144] = 16'b0000000011100011;
    cells[145] = 16'b0000000011100001;
    cells[146] = 16'b0000000011100000;
    cells[147] = 16'b0000000011011110;
    cells[148] = 16'b0000000011011101;
    cells[149] = 16'b0000000011011011;
    cells[150] = 16'b0000000011011010;
    cells[151] = 16'b0000000011011001;
    cells[152] = 16'b0000000011010111;
    cells[153] = 16'b0000000011010110;
    cells[154] = 16'b0000000011010100;
    cells[155] = 16'b0000000011010011;
    cells[156] = 16'b0000000011010010;
    cells[157] = 16'b0000000011010000;
    cells[158] = 16'b0000000011001111;
    cells[159] = 16'b0000000011001110;
    cells[160] = 16'b0000000011001100;
    cells[161] = 16'b0000000011001011;
    cells[162] = 16'b0000000011001010;
    cells[163] = 16'b0000000011001001;
    cells[164] = 16'b0000000011000111;
    cells[165] = 16'b0000000011000110;
    cells[166] = 16'b0000000011000101;
    cells[167] = 16'b0000000011000100;
    cells[168] = 16'b0000000011000011;
    cells[169] = 16'b0000000011000001;
    cells[170] = 16'b0000000011000000;
    cells[171] = 16'b0000000010111111;
    cells[172] = 16'b0000000010111110;
    cells[173] = 16'b0000000010111101;
    cells[174] = 16'b0000000010111100;
    cells[175] = 16'b0000000010111011;
    cells[176] = 16'b0000000010111010;
    cells[177] = 16'b0000000010111001;
    cells[178] = 16'b0000000010111000;
    cells[179] = 16'b0000000010110111;
    cells[180] = 16'b0000000010110110;
    cells[181] = 16'b0000000010110101;
    cells[182] = 16'b0000000010110100;
    cells[183] = 16'b0000000010110011;
    cells[184] = 16'b0000000010110010;
    cells[185] = 16'b0000000010110001;
    cells[186] = 16'b0000000010110000;
    cells[187] = 16'b0000000010101111;
    cells[188] = 16'b0000000010101110;
    cells[189] = 16'b0000000010101101;
    cells[190] = 16'b0000000010101100;
    cells[191] = 16'b0000000010101011;
    cells[192] = 16'b0000000010101010;
    cells[193] = 16'b0000000010101001;
    cells[194] = 16'b0000000010101000;
    cells[195] = 16'b0000000010101000;
    cells[196] = 16'b0000000010100111;
    cells[197] = 16'b0000000010100110;
    cells[198] = 16'b0000000010100101;
    cells[199] = 16'b0000000010100100;
    cells[200] = 16'b0000000010100011;
    cells[201] = 16'b0000000010100011;
    cells[202] = 16'b0000000010100010;
    cells[203] = 16'b0000000010100001;
    cells[204] = 16'b0000000010100000;
    cells[205] = 16'b0000000010011111;
    cells[206] = 16'b0000000010011111;
    cells[207] = 16'b0000000010011110;
    cells[208] = 16'b0000000010011101;
    cells[209] = 16'b0000000010011100;
    cells[210] = 16'b0000000010011100;
    cells[211] = 16'b0000000010011011;
    cells[212] = 16'b0000000010011010;
    cells[213] = 16'b0000000010011001;
    cells[214] = 16'b0000000010011001;
    cells[215] = 16'b0000000010011000;
    cells[216] = 16'b0000000010010111;
    cells[217] = 16'b0000000010010111;
    cells[218] = 16'b0000000010010110;
    cells[219] = 16'b0000000010010101;
    cells[220] = 16'b0000000010010100;
    cells[221] = 16'b0000000010010100;
    cells[222] = 16'b0000000010010011;
    cells[223] = 16'b0000000010010010;
    cells[224] = 16'b0000000010010010;
    cells[225] = 16'b0000000010010001;
    cells[226] = 16'b0000000010010000;
    cells[227] = 16'b0000000010010000;
    cells[228] = 16'b0000000010001111;
    cells[229] = 16'b0000000010001111;
    cells[230] = 16'b0000000010001110;
    cells[231] = 16'b0000000010001101;
    cells[232] = 16'b0000000010001101;
    cells[233] = 16'b0000000010001100;
    cells[234] = 16'b0000000010001100;
    cells[235] = 16'b0000000010001011;
    cells[236] = 16'b0000000010001010;
    cells[237] = 16'b0000000010001010;
    cells[238] = 16'b0000000010001001;
    cells[239] = 16'b0000000010001001;
    cells[240] = 16'b0000000010001000;
    cells[241] = 16'b0000000010000111;
    cells[242] = 16'b0000000010000111;
    cells[243] = 16'b0000000010000110;
    cells[244] = 16'b0000000010000110;
    cells[245] = 16'b0000000010000101;
    cells[246] = 16'b0000000010000101;
    cells[247] = 16'b0000000010000100;
    cells[248] = 16'b0000000010000100;
    cells[249] = 16'b0000000010000011;
    cells[250] = 16'b0000000010000011;
    cells[251] = 16'b0000000010000010;
    cells[252] = 16'b0000000010000010;
    cells[253] = 16'b0000000010000001;
    cells[254] = 16'b0000000010000001;
    cells[255] = 16'b0000000010000000;
    cells[256] = 16'b0000000010000000;
    cells[257] = 16'b0000000001111111;
    cells[258] = 16'b0000000001111111;
    cells[259] = 16'b0000000001111110;
    cells[260] = 16'b0000000001111110;
    cells[261] = 16'b0000000001111101;
    cells[262] = 16'b0000000001111101;
    cells[263] = 16'b0000000001111100;
    cells[264] = 16'b0000000001111100;
    cells[265] = 16'b0000000001111011;
    cells[266] = 16'b0000000001111011;
    cells[267] = 16'b0000000001111010;
    cells[268] = 16'b0000000001111010;
    cells[269] = 16'b0000000001111001;
    cells[270] = 16'b0000000001111001;
    cells[271] = 16'b0000000001111000;
    cells[272] = 16'b0000000001111000;
    cells[273] = 16'b0000000001111000;
    cells[274] = 16'b0000000001110111;
    cells[275] = 16'b0000000001110111;
    cells[276] = 16'b0000000001110110;
    cells[277] = 16'b0000000001110110;
    cells[278] = 16'b0000000001110101;
    cells[279] = 16'b0000000001110101;
    cells[280] = 16'b0000000001110101;
    cells[281] = 16'b0000000001110100;
    cells[282] = 16'b0000000001110100;
    cells[283] = 16'b0000000001110011;
    cells[284] = 16'b0000000001110011;
    cells[285] = 16'b0000000001110010;
    cells[286] = 16'b0000000001110010;
    cells[287] = 16'b0000000001110010;
    cells[288] = 16'b0000000001110001;
    cells[289] = 16'b0000000001110001;
    cells[290] = 16'b0000000001110000;
    cells[291] = 16'b0000000001110000;
    cells[292] = 16'b0000000001110000;
    cells[293] = 16'b0000000001101111;
    cells[294] = 16'b0000000001101111;
    cells[295] = 16'b0000000001101111;
    cells[296] = 16'b0000000001101110;
    cells[297] = 16'b0000000001101110;
    cells[298] = 16'b0000000001101101;
    cells[299] = 16'b0000000001101101;
    cells[300] = 16'b0000000001101101;
    cells[301] = 16'b0000000001101100;
    cells[302] = 16'b0000000001101100;
    cells[303] = 16'b0000000001101100;
    cells[304] = 16'b0000000001101011;
    cells[305] = 16'b0000000001101011;
    cells[306] = 16'b0000000001101011;
    cells[307] = 16'b0000000001101010;
    cells[308] = 16'b0000000001101010;
    cells[309] = 16'b0000000001101010;
    cells[310] = 16'b0000000001101001;
    cells[311] = 16'b0000000001101001;
    cells[312] = 16'b0000000001101001;
    cells[313] = 16'b0000000001101000;
    cells[314] = 16'b0000000001101000;
    cells[315] = 16'b0000000001101000;
    cells[316] = 16'b0000000001100111;
    cells[317] = 16'b0000000001100111;
    cells[318] = 16'b0000000001100111;
    cells[319] = 16'b0000000001100110;
    cells[320] = 16'b0000000001100110;
    cells[321] = 16'b0000000001100110;
    cells[322] = 16'b0000000001100101;
    cells[323] = 16'b0000000001100101;
    cells[324] = 16'b0000000001100101;
    cells[325] = 16'b0000000001100100;
    cells[326] = 16'b0000000001100100;
    cells[327] = 16'b0000000001100100;
    cells[328] = 16'b0000000001100011;
    cells[329] = 16'b0000000001100011;
    cells[330] = 16'b0000000001100011;
    cells[331] = 16'b0000000001100010;
    cells[332] = 16'b0000000001100010;
    cells[333] = 16'b0000000001100010;
    cells[334] = 16'b0000000001100010;
    cells[335] = 16'b0000000001100001;
    cells[336] = 16'b0000000001100001;
    cells[337] = 16'b0000000001100001;
    cells[338] = 16'b0000000001100000;
    cells[339] = 16'b0000000001100000;
    cells[340] = 16'b0000000001100000;
    cells[341] = 16'b0000000001100000;
    cells[342] = 16'b0000000001011111;
    cells[343] = 16'b0000000001011111;
    cells[344] = 16'b0000000001011111;
    cells[345] = 16'b0000000001011110;
    cells[346] = 16'b0000000001011110;
    cells[347] = 16'b0000000001011110;
    cells[348] = 16'b0000000001011110;
    cells[349] = 16'b0000000001011101;
    cells[350] = 16'b0000000001011101;
    cells[351] = 16'b0000000001011101;
    cells[352] = 16'b0000000001011101;
    cells[353] = 16'b0000000001011100;
    cells[354] = 16'b0000000001011100;
    cells[355] = 16'b0000000001011100;
    cells[356] = 16'b0000000001011100;
    cells[357] = 16'b0000000001011011;
    cells[358] = 16'b0000000001011011;
    cells[359] = 16'b0000000001011011;
    cells[360] = 16'b0000000001011011;
    cells[361] = 16'b0000000001011010;
    cells[362] = 16'b0000000001011010;
    cells[363] = 16'b0000000001011010;
    cells[364] = 16'b0000000001011010;
    cells[365] = 16'b0000000001011001;
    cells[366] = 16'b0000000001011001;
    cells[367] = 16'b0000000001011001;
    cells[368] = 16'b0000000001011001;
    cells[369] = 16'b0000000001011000;
    cells[370] = 16'b0000000001011000;
    cells[371] = 16'b0000000001011000;
    cells[372] = 16'b0000000001011000;
    cells[373] = 16'b0000000001010111;
    cells[374] = 16'b0000000001010111;
    cells[375] = 16'b0000000001010111;
    cells[376] = 16'b0000000001010111;
    cells[377] = 16'b0000000001010110;
    cells[378] = 16'b0000000001010110;
    cells[379] = 16'b0000000001010110;
    cells[380] = 16'b0000000001010110;
    cells[381] = 16'b0000000001010110;
    cells[382] = 16'b0000000001010101;
    cells[383] = 16'b0000000001010101;
    cells[384] = 16'b0000000001010101;
    cells[385] = 16'b0000000001010101;
    cells[386] = 16'b0000000001010100;
    cells[387] = 16'b0000000001010100;
    cells[388] = 16'b0000000001010100;
    cells[389] = 16'b0000000001010100;
    cells[390] = 16'b0000000001010100;
    cells[391] = 16'b0000000001010011;
    cells[392] = 16'b0000000001010011;
    cells[393] = 16'b0000000001010011;
    cells[394] = 16'b0000000001010011;
    cells[395] = 16'b0000000001010010;
    cells[396] = 16'b0000000001010010;
    cells[397] = 16'b0000000001010010;
    cells[398] = 16'b0000000001010010;
    cells[399] = 16'b0000000001010010;
    cells[400] = 16'b0000000001010001;
    cells[401] = 16'b0000000001010001;
    cells[402] = 16'b0000000001010001;
    cells[403] = 16'b0000000001010001;
    cells[404] = 16'b0000000001010001;
    cells[405] = 16'b0000000001010000;
    cells[406] = 16'b0000000001010000;
    cells[407] = 16'b0000000001010000;
    cells[408] = 16'b0000000001010000;
    cells[409] = 16'b0000000001010000;
    cells[410] = 16'b0000000001001111;
    cells[411] = 16'b0000000001001111;
    cells[412] = 16'b0000000001001111;
    cells[413] = 16'b0000000001001111;
    cells[414] = 16'b0000000001001111;
    cells[415] = 16'b0000000001001110;
    cells[416] = 16'b0000000001001110;
    cells[417] = 16'b0000000001001110;
    cells[418] = 16'b0000000001001110;
    cells[419] = 16'b0000000001001110;
    cells[420] = 16'b0000000001001110;
    cells[421] = 16'b0000000001001101;
    cells[422] = 16'b0000000001001101;
    cells[423] = 16'b0000000001001101;
    cells[424] = 16'b0000000001001101;
    cells[425] = 16'b0000000001001101;
    cells[426] = 16'b0000000001001100;
    cells[427] = 16'b0000000001001100;
    cells[428] = 16'b0000000001001100;
    cells[429] = 16'b0000000001001100;
    cells[430] = 16'b0000000001001100;
    cells[431] = 16'b0000000001001100;
    cells[432] = 16'b0000000001001011;
    cells[433] = 16'b0000000001001011;
    cells[434] = 16'b0000000001001011;
    cells[435] = 16'b0000000001001011;
    cells[436] = 16'b0000000001001011;
    cells[437] = 16'b0000000001001010;
    cells[438] = 16'b0000000001001010;
    cells[439] = 16'b0000000001001010;
    cells[440] = 16'b0000000001001010;
    cells[441] = 16'b0000000001001010;
    cells[442] = 16'b0000000001001010;
    cells[443] = 16'b0000000001001001;
    cells[444] = 16'b0000000001001001;
    cells[445] = 16'b0000000001001001;
    cells[446] = 16'b0000000001001001;
    cells[447] = 16'b0000000001001001;
    cells[448] = 16'b0000000001001001;
    cells[449] = 16'b0000000001001000;
    cells[450] = 16'b0000000001001000;
    cells[451] = 16'b0000000001001000;
    cells[452] = 16'b0000000001001000;
    cells[453] = 16'b0000000001001000;
    cells[454] = 16'b0000000001001000;
    cells[455] = 16'b0000000001001000;
    cells[456] = 16'b0000000001000111;
    cells[457] = 16'b0000000001000111;
    cells[458] = 16'b0000000001000111;
    cells[459] = 16'b0000000001000111;
    cells[460] = 16'b0000000001000111;
    cells[461] = 16'b0000000001000111;
    cells[462] = 16'b0000000001000110;
    cells[463] = 16'b0000000001000110;
    cells[464] = 16'b0000000001000110;
    cells[465] = 16'b0000000001000110;
    cells[466] = 16'b0000000001000110;
    cells[467] = 16'b0000000001000110;
    cells[468] = 16'b0000000001000110;
    cells[469] = 16'b0000000001000101;
    cells[470] = 16'b0000000001000101;
    cells[471] = 16'b0000000001000101;
    cells[472] = 16'b0000000001000101;
    cells[473] = 16'b0000000001000101;
    cells[474] = 16'b0000000001000101;
    cells[475] = 16'b0000000001000100;
    cells[476] = 16'b0000000001000100;
    cells[477] = 16'b0000000001000100;
    cells[478] = 16'b0000000001000100;
    cells[479] = 16'b0000000001000100;
    cells[480] = 16'b0000000001000100;
    cells[481] = 16'b0000000001000100;
    cells[482] = 16'b0000000001000011;
    cells[483] = 16'b0000000001000011;
    cells[484] = 16'b0000000001000011;
    cells[485] = 16'b0000000001000011;
    cells[486] = 16'b0000000001000011;
    cells[487] = 16'b0000000001000011;
    cells[488] = 16'b0000000001000011;
    cells[489] = 16'b0000000001000011;
    cells[490] = 16'b0000000001000010;
    cells[491] = 16'b0000000001000010;
    cells[492] = 16'b0000000001000010;
    cells[493] = 16'b0000000001000010;
    cells[494] = 16'b0000000001000010;
    cells[495] = 16'b0000000001000010;
    cells[496] = 16'b0000000001000010;
    cells[497] = 16'b0000000001000001;
    cells[498] = 16'b0000000001000001;
    cells[499] = 16'b0000000001000001;
    cells[500] = 16'b0000000001000001;
    cells[501] = 16'b0000000001000001;
    cells[502] = 16'b0000000001000001;
    cells[503] = 16'b0000000001000001;
    cells[504] = 16'b0000000001000001;
    cells[505] = 16'b0000000001000000;
    cells[506] = 16'b0000000001000000;
    cells[507] = 16'b0000000001000000;
    cells[508] = 16'b0000000001000000;
    cells[509] = 16'b0000000001000000;
    cells[510] = 16'b0000000001000000;
    cells[511] = 16'b0000000001000000;
    cells[512] = 16'b0000000001000000;
    cells[513] = 16'b0000000000111111;
    cells[514] = 16'b0000000000111111;
    cells[515] = 16'b0000000000111111;
    cells[516] = 16'b0000000000111111;
    cells[517] = 16'b0000000000111111;
    cells[518] = 16'b0000000000111111;
    cells[519] = 16'b0000000000111111;
    cells[520] = 16'b0000000000111111;
    cells[521] = 16'b0000000000111110;
    cells[522] = 16'b0000000000111110;
    cells[523] = 16'b0000000000111110;
    cells[524] = 16'b0000000000111110;
    cells[525] = 16'b0000000000111110;
    cells[526] = 16'b0000000000111110;
    cells[527] = 16'b0000000000111110;
    cells[528] = 16'b0000000000111110;
    cells[529] = 16'b0000000000111101;
    cells[530] = 16'b0000000000111101;
    cells[531] = 16'b0000000000111101;
    cells[532] = 16'b0000000000111101;
    cells[533] = 16'b0000000000111101;
    cells[534] = 16'b0000000000111101;
    cells[535] = 16'b0000000000111101;
    cells[536] = 16'b0000000000111101;
    cells[537] = 16'b0000000000111101;
    cells[538] = 16'b0000000000111100;
    cells[539] = 16'b0000000000111100;
    cells[540] = 16'b0000000000111100;
    cells[541] = 16'b0000000000111100;
    cells[542] = 16'b0000000000111100;
    cells[543] = 16'b0000000000111100;
    cells[544] = 16'b0000000000111100;
    cells[545] = 16'b0000000000111100;
    cells[546] = 16'b0000000000111100;
    cells[547] = 16'b0000000000111011;
    cells[548] = 16'b0000000000111011;
    cells[549] = 16'b0000000000111011;
    cells[550] = 16'b0000000000111011;
    cells[551] = 16'b0000000000111011;
    cells[552] = 16'b0000000000111011;
    cells[553] = 16'b0000000000111011;
    cells[554] = 16'b0000000000111011;
    cells[555] = 16'b0000000000111011;
    cells[556] = 16'b0000000000111010;
    cells[557] = 16'b0000000000111010;
    cells[558] = 16'b0000000000111010;
    cells[559] = 16'b0000000000111010;
    cells[560] = 16'b0000000000111010;
    cells[561] = 16'b0000000000111010;
    cells[562] = 16'b0000000000111010;
    cells[563] = 16'b0000000000111010;
    cells[564] = 16'b0000000000111010;
    cells[565] = 16'b0000000000111001;
    cells[566] = 16'b0000000000111001;
    cells[567] = 16'b0000000000111001;
    cells[568] = 16'b0000000000111001;
    cells[569] = 16'b0000000000111001;
    cells[570] = 16'b0000000000111001;
    cells[571] = 16'b0000000000111001;
    cells[572] = 16'b0000000000111001;
    cells[573] = 16'b0000000000111001;
    cells[574] = 16'b0000000000111001;
    cells[575] = 16'b0000000000111000;
    cells[576] = 16'b0000000000111000;
    cells[577] = 16'b0000000000111000;
    cells[578] = 16'b0000000000111000;
    cells[579] = 16'b0000000000111000;
    cells[580] = 16'b0000000000111000;
    cells[581] = 16'b0000000000111000;
    cells[582] = 16'b0000000000111000;
    cells[583] = 16'b0000000000111000;
    cells[584] = 16'b0000000000111000;
    cells[585] = 16'b0000000000111000;
    cells[586] = 16'b0000000000110111;
    cells[587] = 16'b0000000000110111;
    cells[588] = 16'b0000000000110111;
    cells[589] = 16'b0000000000110111;
    cells[590] = 16'b0000000000110111;
    cells[591] = 16'b0000000000110111;
    cells[592] = 16'b0000000000110111;
    cells[593] = 16'b0000000000110111;
    cells[594] = 16'b0000000000110111;
    cells[595] = 16'b0000000000110111;
    cells[596] = 16'b0000000000110110;
    cells[597] = 16'b0000000000110110;
    cells[598] = 16'b0000000000110110;
    cells[599] = 16'b0000000000110110;
    cells[600] = 16'b0000000000110110;
    cells[601] = 16'b0000000000110110;
    cells[602] = 16'b0000000000110110;
    cells[603] = 16'b0000000000110110;
    cells[604] = 16'b0000000000110110;
    cells[605] = 16'b0000000000110110;
    cells[606] = 16'b0000000000110110;
    cells[607] = 16'b0000000000110101;
    cells[608] = 16'b0000000000110101;
    cells[609] = 16'b0000000000110101;
    cells[610] = 16'b0000000000110101;
    cells[611] = 16'b0000000000110101;
    cells[612] = 16'b0000000000110101;
    cells[613] = 16'b0000000000110101;
    cells[614] = 16'b0000000000110101;
    cells[615] = 16'b0000000000110101;
    cells[616] = 16'b0000000000110101;
    cells[617] = 16'b0000000000110101;
    cells[618] = 16'b0000000000110101;
    cells[619] = 16'b0000000000110100;
    cells[620] = 16'b0000000000110100;
    cells[621] = 16'b0000000000110100;
    cells[622] = 16'b0000000000110100;
    cells[623] = 16'b0000000000110100;
    cells[624] = 16'b0000000000110100;
    cells[625] = 16'b0000000000110100;
    cells[626] = 16'b0000000000110100;
    cells[627] = 16'b0000000000110100;
    cells[628] = 16'b0000000000110100;
    cells[629] = 16'b0000000000110100;
    cells[630] = 16'b0000000000110100;
    cells[631] = 16'b0000000000110011;
    cells[632] = 16'b0000000000110011;
    cells[633] = 16'b0000000000110011;
    cells[634] = 16'b0000000000110011;
    cells[635] = 16'b0000000000110011;
    cells[636] = 16'b0000000000110011;
    cells[637] = 16'b0000000000110011;
    cells[638] = 16'b0000000000110011;
    cells[639] = 16'b0000000000110011;
    cells[640] = 16'b0000000000110011;
    cells[641] = 16'b0000000000110011;
    cells[642] = 16'b0000000000110011;
    cells[643] = 16'b0000000000110010;
    cells[644] = 16'b0000000000110010;
    cells[645] = 16'b0000000000110010;
    cells[646] = 16'b0000000000110010;
    cells[647] = 16'b0000000000110010;
    cells[648] = 16'b0000000000110010;
    cells[649] = 16'b0000000000110010;
    cells[650] = 16'b0000000000110010;
    cells[651] = 16'b0000000000110010;
    cells[652] = 16'b0000000000110010;
    cells[653] = 16'b0000000000110010;
    cells[654] = 16'b0000000000110010;
    cells[655] = 16'b0000000000110010;
    cells[656] = 16'b0000000000110001;
    cells[657] = 16'b0000000000110001;
    cells[658] = 16'b0000000000110001;
    cells[659] = 16'b0000000000110001;
    cells[660] = 16'b0000000000110001;
    cells[661] = 16'b0000000000110001;
    cells[662] = 16'b0000000000110001;
    cells[663] = 16'b0000000000110001;
    cells[664] = 16'b0000000000110001;
    cells[665] = 16'b0000000000110001;
    cells[666] = 16'b0000000000110001;
    cells[667] = 16'b0000000000110001;
    cells[668] = 16'b0000000000110001;
    cells[669] = 16'b0000000000110000;
    cells[670] = 16'b0000000000110000;
    cells[671] = 16'b0000000000110000;
    cells[672] = 16'b0000000000110000;
    cells[673] = 16'b0000000000110000;
    cells[674] = 16'b0000000000110000;
    cells[675] = 16'b0000000000110000;
    cells[676] = 16'b0000000000110000;
    cells[677] = 16'b0000000000110000;
    cells[678] = 16'b0000000000110000;
    cells[679] = 16'b0000000000110000;
    cells[680] = 16'b0000000000110000;
    cells[681] = 16'b0000000000110000;
    cells[682] = 16'b0000000000110000;
    cells[683] = 16'b0000000000101111;
    cells[684] = 16'b0000000000101111;
    cells[685] = 16'b0000000000101111;
    cells[686] = 16'b0000000000101111;
    cells[687] = 16'b0000000000101111;
    cells[688] = 16'b0000000000101111;
    cells[689] = 16'b0000000000101111;
    cells[690] = 16'b0000000000101111;
    cells[691] = 16'b0000000000101111;
    cells[692] = 16'b0000000000101111;
    cells[693] = 16'b0000000000101111;
    cells[694] = 16'b0000000000101111;
    cells[695] = 16'b0000000000101111;
    cells[696] = 16'b0000000000101111;
    cells[697] = 16'b0000000000101111;
    cells[698] = 16'b0000000000101110;
    cells[699] = 16'b0000000000101110;
    cells[700] = 16'b0000000000101110;
    cells[701] = 16'b0000000000101110;
    cells[702] = 16'b0000000000101110;
    cells[703] = 16'b0000000000101110;
    cells[704] = 16'b0000000000101110;
    cells[705] = 16'b0000000000101110;
    cells[706] = 16'b0000000000101110;
    cells[707] = 16'b0000000000101110;
    cells[708] = 16'b0000000000101110;
    cells[709] = 16'b0000000000101110;
    cells[710] = 16'b0000000000101110;
    cells[711] = 16'b0000000000101110;
    cells[712] = 16'b0000000000101110;
    cells[713] = 16'b0000000000101101;
    cells[714] = 16'b0000000000101101;
    cells[715] = 16'b0000000000101101;
    cells[716] = 16'b0000000000101101;
    cells[717] = 16'b0000000000101101;
    cells[718] = 16'b0000000000101101;
    cells[719] = 16'b0000000000101101;
    cells[720] = 16'b0000000000101101;
    cells[721] = 16'b0000000000101101;
    cells[722] = 16'b0000000000101101;
    cells[723] = 16'b0000000000101101;
    cells[724] = 16'b0000000000101101;
    cells[725] = 16'b0000000000101101;
    cells[726] = 16'b0000000000101101;
    cells[727] = 16'b0000000000101101;
    cells[728] = 16'b0000000000101101;
    cells[729] = 16'b0000000000101100;
    cells[730] = 16'b0000000000101100;
    cells[731] = 16'b0000000000101100;
    cells[732] = 16'b0000000000101100;
    cells[733] = 16'b0000000000101100;
    cells[734] = 16'b0000000000101100;
    cells[735] = 16'b0000000000101100;
    cells[736] = 16'b0000000000101100;
    cells[737] = 16'b0000000000101100;
    cells[738] = 16'b0000000000101100;
    cells[739] = 16'b0000000000101100;
    cells[740] = 16'b0000000000101100;
    cells[741] = 16'b0000000000101100;
    cells[742] = 16'b0000000000101100;
    cells[743] = 16'b0000000000101100;
    cells[744] = 16'b0000000000101100;
    cells[745] = 16'b0000000000101011;
    cells[746] = 16'b0000000000101011;
    cells[747] = 16'b0000000000101011;
    cells[748] = 16'b0000000000101011;
    cells[749] = 16'b0000000000101011;
    cells[750] = 16'b0000000000101011;
    cells[751] = 16'b0000000000101011;
    cells[752] = 16'b0000000000101011;
    cells[753] = 16'b0000000000101011;
    cells[754] = 16'b0000000000101011;
    cells[755] = 16'b0000000000101011;
    cells[756] = 16'b0000000000101011;
    cells[757] = 16'b0000000000101011;
    cells[758] = 16'b0000000000101011;
    cells[759] = 16'b0000000000101011;
    cells[760] = 16'b0000000000101011;
    cells[761] = 16'b0000000000101011;
    cells[762] = 16'b0000000000101011;
    cells[763] = 16'b0000000000101010;
    cells[764] = 16'b0000000000101010;
    cells[765] = 16'b0000000000101010;
    cells[766] = 16'b0000000000101010;
    cells[767] = 16'b0000000000101010;
    cells[768] = 16'b0000000000101010;
    cells[769] = 16'b0000000000101010;
    cells[770] = 16'b0000000000101010;
    cells[771] = 16'b0000000000101010;
    cells[772] = 16'b0000000000101010;
    cells[773] = 16'b0000000000101010;
    cells[774] = 16'b0000000000101010;
    cells[775] = 16'b0000000000101010;
    cells[776] = 16'b0000000000101010;
    cells[777] = 16'b0000000000101010;
    cells[778] = 16'b0000000000101010;
    cells[779] = 16'b0000000000101010;
    cells[780] = 16'b0000000000101010;
    cells[781] = 16'b0000000000101001;
    cells[782] = 16'b0000000000101001;
    cells[783] = 16'b0000000000101001;
    cells[784] = 16'b0000000000101001;
    cells[785] = 16'b0000000000101001;
    cells[786] = 16'b0000000000101001;
    cells[787] = 16'b0000000000101001;
    cells[788] = 16'b0000000000101001;
    cells[789] = 16'b0000000000101001;
    cells[790] = 16'b0000000000101001;
    cells[791] = 16'b0000000000101001;
    cells[792] = 16'b0000000000101001;
    cells[793] = 16'b0000000000101001;
    cells[794] = 16'b0000000000101001;
    cells[795] = 16'b0000000000101001;
    cells[796] = 16'b0000000000101001;
    cells[797] = 16'b0000000000101001;
    cells[798] = 16'b0000000000101001;
    cells[799] = 16'b0000000000101001;
    cells[800] = 16'b0000000000101000;
    cells[801] = 16'b0000000000101000;
    cells[802] = 16'b0000000000101000;
    cells[803] = 16'b0000000000101000;
    cells[804] = 16'b0000000000101000;
    cells[805] = 16'b0000000000101000;
    cells[806] = 16'b0000000000101000;
    cells[807] = 16'b0000000000101000;
    cells[808] = 16'b0000000000101000;
    cells[809] = 16'b0000000000101000;
    cells[810] = 16'b0000000000101000;
    cells[811] = 16'b0000000000101000;
    cells[812] = 16'b0000000000101000;
    cells[813] = 16'b0000000000101000;
    cells[814] = 16'b0000000000101000;
    cells[815] = 16'b0000000000101000;
    cells[816] = 16'b0000000000101000;
    cells[817] = 16'b0000000000101000;
    cells[818] = 16'b0000000000101000;
    cells[819] = 16'b0000000000101000;
    cells[820] = 16'b0000000000100111;
    cells[821] = 16'b0000000000100111;
    cells[822] = 16'b0000000000100111;
    cells[823] = 16'b0000000000100111;
    cells[824] = 16'b0000000000100111;
    cells[825] = 16'b0000000000100111;
    cells[826] = 16'b0000000000100111;
    cells[827] = 16'b0000000000100111;
    cells[828] = 16'b0000000000100111;
    cells[829] = 16'b0000000000100111;
    cells[830] = 16'b0000000000100111;
    cells[831] = 16'b0000000000100111;
    cells[832] = 16'b0000000000100111;
    cells[833] = 16'b0000000000100111;
    cells[834] = 16'b0000000000100111;
    cells[835] = 16'b0000000000100111;
    cells[836] = 16'b0000000000100111;
    cells[837] = 16'b0000000000100111;
    cells[838] = 16'b0000000000100111;
    cells[839] = 16'b0000000000100111;
    cells[840] = 16'b0000000000100111;
    cells[841] = 16'b0000000000100110;
    cells[842] = 16'b0000000000100110;
    cells[843] = 16'b0000000000100110;
    cells[844] = 16'b0000000000100110;
    cells[845] = 16'b0000000000100110;
    cells[846] = 16'b0000000000100110;
    cells[847] = 16'b0000000000100110;
    cells[848] = 16'b0000000000100110;
    cells[849] = 16'b0000000000100110;
    cells[850] = 16'b0000000000100110;
    cells[851] = 16'b0000000000100110;
    cells[852] = 16'b0000000000100110;
    cells[853] = 16'b0000000000100110;
    cells[854] = 16'b0000000000100110;
    cells[855] = 16'b0000000000100110;
    cells[856] = 16'b0000000000100110;
    cells[857] = 16'b0000000000100110;
    cells[858] = 16'b0000000000100110;
    cells[859] = 16'b0000000000100110;
    cells[860] = 16'b0000000000100110;
    cells[861] = 16'b0000000000100110;
    cells[862] = 16'b0000000000100110;
    cells[863] = 16'b0000000000100101;
    cells[864] = 16'b0000000000100101;
    cells[865] = 16'b0000000000100101;
    cells[866] = 16'b0000000000100101;
    cells[867] = 16'b0000000000100101;
    cells[868] = 16'b0000000000100101;
    cells[869] = 16'b0000000000100101;
    cells[870] = 16'b0000000000100101;
    cells[871] = 16'b0000000000100101;
    cells[872] = 16'b0000000000100101;
    cells[873] = 16'b0000000000100101;
    cells[874] = 16'b0000000000100101;
    cells[875] = 16'b0000000000100101;
    cells[876] = 16'b0000000000100101;
    cells[877] = 16'b0000000000100101;
    cells[878] = 16'b0000000000100101;
    cells[879] = 16'b0000000000100101;
    cells[880] = 16'b0000000000100101;
    cells[881] = 16'b0000000000100101;
    cells[882] = 16'b0000000000100101;
    cells[883] = 16'b0000000000100101;
    cells[884] = 16'b0000000000100101;
    cells[885] = 16'b0000000000100101;
    cells[886] = 16'b0000000000100100;
    cells[887] = 16'b0000000000100100;
    cells[888] = 16'b0000000000100100;
    cells[889] = 16'b0000000000100100;
    cells[890] = 16'b0000000000100100;
    cells[891] = 16'b0000000000100100;
    cells[892] = 16'b0000000000100100;
    cells[893] = 16'b0000000000100100;
    cells[894] = 16'b0000000000100100;
    cells[895] = 16'b0000000000100100;
    cells[896] = 16'b0000000000100100;
    cells[897] = 16'b0000000000100100;
    cells[898] = 16'b0000000000100100;
    cells[899] = 16'b0000000000100100;
    cells[900] = 16'b0000000000100100;
    cells[901] = 16'b0000000000100100;
    cells[902] = 16'b0000000000100100;
    cells[903] = 16'b0000000000100100;
    cells[904] = 16'b0000000000100100;
    cells[905] = 16'b0000000000100100;
    cells[906] = 16'b0000000000100100;
    cells[907] = 16'b0000000000100100;
    cells[908] = 16'b0000000000100100;
    cells[909] = 16'b0000000000100100;
    cells[910] = 16'b0000000000100100;
    cells[911] = 16'b0000000000100011;
    cells[912] = 16'b0000000000100011;
    cells[913] = 16'b0000000000100011;
    cells[914] = 16'b0000000000100011;
    cells[915] = 16'b0000000000100011;
    cells[916] = 16'b0000000000100011;
    cells[917] = 16'b0000000000100011;
    cells[918] = 16'b0000000000100011;
    cells[919] = 16'b0000000000100011;
    cells[920] = 16'b0000000000100011;
    cells[921] = 16'b0000000000100011;
    cells[922] = 16'b0000000000100011;
    cells[923] = 16'b0000000000100011;
    cells[924] = 16'b0000000000100011;
    cells[925] = 16'b0000000000100011;
    cells[926] = 16'b0000000000100011;
    cells[927] = 16'b0000000000100011;
    cells[928] = 16'b0000000000100011;
    cells[929] = 16'b0000000000100011;
    cells[930] = 16'b0000000000100011;
    cells[931] = 16'b0000000000100011;
    cells[932] = 16'b0000000000100011;
    cells[933] = 16'b0000000000100011;
    cells[934] = 16'b0000000000100011;
    cells[935] = 16'b0000000000100011;
    cells[936] = 16'b0000000000100011;
    cells[937] = 16'b0000000000100010;
    cells[938] = 16'b0000000000100010;
    cells[939] = 16'b0000000000100010;
    cells[940] = 16'b0000000000100010;
    cells[941] = 16'b0000000000100010;
    cells[942] = 16'b0000000000100010;
    cells[943] = 16'b0000000000100010;
    cells[944] = 16'b0000000000100010;
    cells[945] = 16'b0000000000100010;
    cells[946] = 16'b0000000000100010;
    cells[947] = 16'b0000000000100010;
    cells[948] = 16'b0000000000100010;
    cells[949] = 16'b0000000000100010;
    cells[950] = 16'b0000000000100010;
    cells[951] = 16'b0000000000100010;
    cells[952] = 16'b0000000000100010;
    cells[953] = 16'b0000000000100010;
    cells[954] = 16'b0000000000100010;
    cells[955] = 16'b0000000000100010;
    cells[956] = 16'b0000000000100010;
    cells[957] = 16'b0000000000100010;
    cells[958] = 16'b0000000000100010;
    cells[959] = 16'b0000000000100010;
    cells[960] = 16'b0000000000100010;
    cells[961] = 16'b0000000000100010;
    cells[962] = 16'b0000000000100010;
    cells[963] = 16'b0000000000100010;
    cells[964] = 16'b0000000000100001;
    cells[965] = 16'b0000000000100001;
    cells[966] = 16'b0000000000100001;
    cells[967] = 16'b0000000000100001;
    cells[968] = 16'b0000000000100001;
    cells[969] = 16'b0000000000100001;
    cells[970] = 16'b0000000000100001;
    cells[971] = 16'b0000000000100001;
    cells[972] = 16'b0000000000100001;
    cells[973] = 16'b0000000000100001;
    cells[974] = 16'b0000000000100001;
    cells[975] = 16'b0000000000100001;
    cells[976] = 16'b0000000000100001;
    cells[977] = 16'b0000000000100001;
    cells[978] = 16'b0000000000100001;
    cells[979] = 16'b0000000000100001;
    cells[980] = 16'b0000000000100001;
    cells[981] = 16'b0000000000100001;
    cells[982] = 16'b0000000000100001;
    cells[983] = 16'b0000000000100001;
    cells[984] = 16'b0000000000100001;
    cells[985] = 16'b0000000000100001;
    cells[986] = 16'b0000000000100001;
    cells[987] = 16'b0000000000100001;
    cells[988] = 16'b0000000000100001;
    cells[989] = 16'b0000000000100001;
    cells[990] = 16'b0000000000100001;
    cells[991] = 16'b0000000000100001;
    cells[992] = 16'b0000000000100001;
    cells[993] = 16'b0000000000100000;
    cells[994] = 16'b0000000000100000;
    cells[995] = 16'b0000000000100000;
    cells[996] = 16'b0000000000100000;
    cells[997] = 16'b0000000000100000;
    cells[998] = 16'b0000000000100000;
    cells[999] = 16'b0000000000100000;
    cells[1000] = 16'b0000000000100000;
    cells[1001] = 16'b0000000000100000;
    cells[1002] = 16'b0000000000100000;
    cells[1003] = 16'b0000000000100000;
    cells[1004] = 16'b0000000000100000;
    cells[1005] = 16'b0000000000100000;
    cells[1006] = 16'b0000000000100000;
    cells[1007] = 16'b0000000000100000;
    cells[1008] = 16'b0000000000100000;
    cells[1009] = 16'b0000000000100000;
    cells[1010] = 16'b0000000000100000;
    cells[1011] = 16'b0000000000100000;
    cells[1012] = 16'b0000000000100000;
    cells[1013] = 16'b0000000000100000;
    cells[1014] = 16'b0000000000100000;
    cells[1015] = 16'b0000000000100000;
    cells[1016] = 16'b0000000000100000;
    cells[1017] = 16'b0000000000100000;
    cells[1018] = 16'b0000000000100000;
    cells[1019] = 16'b0000000000100000;
    cells[1020] = 16'b0000000000100000;
    cells[1021] = 16'b0000000000100000;
    cells[1022] = 16'b0000000000100000;
    cells[1023] = 16'b0000000000100000;
end
endmodule

/*Produced by sfl2vl, IP ARCH, Inc. Sun Jul 14 18:45:30 2019
 Licensed to :EVALUATION USER*/
