
/*Produced by sfl2vl, IP ARCH, Inc. Sun Jul 14 18:45:28 2019
 Licensed to :EVALUATION USER*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module sin_table ( p_reset , m_clock , dout , read , angle );
  input p_reset, m_clock;
  wire p_reset, m_clock;
  output [9:0] dout;
  wire [9:0] dout;
  input read;
  wire read;
  input [8:0] angle;
  wire [8:0] angle;
  reg [9:0] dout_reg;
  reg [9:0] cells [0:511];

   assign  dout = dout_reg;
always @(posedge m_clock or posedge p_reset)
  begin
if (p_reset)
     dout_reg <= 10'b0000000000;
else if ((read)) 
      dout_reg <= (cells[angle]);
end
initial begin
    cells[0] = 10'b0000000000;
    cells[1] = 10'b0000000100;
    cells[2] = 10'b0000001000;
    cells[3] = 10'b0000001101;
    cells[4] = 10'b0000010001;
    cells[5] = 10'b0000010110;
    cells[6] = 10'b0000011010;
    cells[7] = 10'b0000011111;
    cells[8] = 10'b0000100011;
    cells[9] = 10'b0000101000;
    cells[10] = 10'b0000101100;
    cells[11] = 10'b0000110000;
    cells[12] = 10'b0000110101;
    cells[13] = 10'b0000111001;
    cells[14] = 10'b0000111101;
    cells[15] = 10'b0001000010;
    cells[16] = 10'b0001000110;
    cells[17] = 10'b0001001010;
    cells[18] = 10'b0001001111;
    cells[19] = 10'b0001010011;
    cells[20] = 10'b0001010111;
    cells[21] = 10'b0001011011;
    cells[22] = 10'b0001011111;
    cells[23] = 10'b0001100100;
    cells[24] = 10'b0001101000;
    cells[25] = 10'b0001101100;
    cells[26] = 10'b0001110000;
    cells[27] = 10'b0001110100;
    cells[28] = 10'b0001111000;
    cells[29] = 10'b0001111100;
    cells[30] = 10'b0010000000;
    cells[31] = 10'b0010000011;
    cells[32] = 10'b0010000111;
    cells[33] = 10'b0010001011;
    cells[34] = 10'b0010001111;
    cells[35] = 10'b0010010010;
    cells[36] = 10'b0010010110;
    cells[37] = 10'b0010011010;
    cells[38] = 10'b0010011101;
    cells[39] = 10'b0010100001;
    cells[40] = 10'b0010100100;
    cells[41] = 10'b0010100111;
    cells[42] = 10'b0010101011;
    cells[43] = 10'b0010101110;
    cells[44] = 10'b0010110001;
    cells[45] = 10'b0010110101;
    cells[46] = 10'b0010111000;
    cells[47] = 10'b0010111011;
    cells[48] = 10'b0010111110;
    cells[49] = 10'b0011000001;
    cells[50] = 10'b0011000100;
    cells[51] = 10'b0011000110;
    cells[52] = 10'b0011001001;
    cells[53] = 10'b0011001100;
    cells[54] = 10'b0011001111;
    cells[55] = 10'b0011010001;
    cells[56] = 10'b0011010100;
    cells[57] = 10'b0011010110;
    cells[58] = 10'b0011011001;
    cells[59] = 10'b0011011011;
    cells[60] = 10'b0011011101;
    cells[61] = 10'b0011011111;
    cells[62] = 10'b0011100010;
    cells[63] = 10'b0011100100;
    cells[64] = 10'b0011100110;
    cells[65] = 10'b0011101000;
    cells[66] = 10'b0011101001;
    cells[67] = 10'b0011101011;
    cells[68] = 10'b0011101101;
    cells[69] = 10'b0011101110;
    cells[70] = 10'b0011110000;
    cells[71] = 10'b0011110010;
    cells[72] = 10'b0011110011;
    cells[73] = 10'b0011110100;
    cells[74] = 10'b0011110110;
    cells[75] = 10'b0011110111;
    cells[76] = 10'b0011111000;
    cells[77] = 10'b0011111001;
    cells[78] = 10'b0011111010;
    cells[79] = 10'b0011111011;
    cells[80] = 10'b0011111100;
    cells[81] = 10'b0011111100;
    cells[82] = 10'b0011111101;
    cells[83] = 10'b0011111110;
    cells[84] = 10'b0011111110;
    cells[85] = 10'b0011111111;
    cells[86] = 10'b0011111111;
    cells[87] = 10'b0011111111;
    cells[88] = 10'b0011111111;
    cells[89] = 10'b0011111111;
    cells[90] = 10'b0100000000;
    cells[91] = 10'b0011111111;
    cells[92] = 10'b0011111111;
    cells[93] = 10'b0011111111;
    cells[94] = 10'b0011111111;
    cells[95] = 10'b0011111111;
    cells[96] = 10'b0011111110;
    cells[97] = 10'b0011111110;
    cells[98] = 10'b0011111101;
    cells[99] = 10'b0011111100;
    cells[100] = 10'b0011111100;
    cells[101] = 10'b0011111011;
    cells[102] = 10'b0011111010;
    cells[103] = 10'b0011111001;
    cells[104] = 10'b0011111000;
    cells[105] = 10'b0011110111;
    cells[106] = 10'b0011110110;
    cells[107] = 10'b0011110100;
    cells[108] = 10'b0011110011;
    cells[109] = 10'b0011110010;
    cells[110] = 10'b0011110000;
    cells[111] = 10'b0011101110;
    cells[112] = 10'b0011101101;
    cells[113] = 10'b0011101011;
    cells[114] = 10'b0011101001;
    cells[115] = 10'b0011101000;
    cells[116] = 10'b0011100110;
    cells[117] = 10'b0011100100;
    cells[118] = 10'b0011100010;
    cells[119] = 10'b0011011111;
    cells[120] = 10'b0011011101;
    cells[121] = 10'b0011011011;
    cells[122] = 10'b0011011001;
    cells[123] = 10'b0011010110;
    cells[124] = 10'b0011010100;
    cells[125] = 10'b0011010001;
    cells[126] = 10'b0011001111;
    cells[127] = 10'b0011001100;
    cells[128] = 10'b0011001001;
    cells[129] = 10'b0011000110;
    cells[130] = 10'b0011000100;
    cells[131] = 10'b0011000001;
    cells[132] = 10'b0010111110;
    cells[133] = 10'b0010111011;
    cells[134] = 10'b0010111000;
    cells[135] = 10'b0010110101;
    cells[136] = 10'b0010110001;
    cells[137] = 10'b0010101110;
    cells[138] = 10'b0010101011;
    cells[139] = 10'b0010100111;
    cells[140] = 10'b0010100100;
    cells[141] = 10'b0010100001;
    cells[142] = 10'b0010011101;
    cells[143] = 10'b0010011010;
    cells[144] = 10'b0010010110;
    cells[145] = 10'b0010010010;
    cells[146] = 10'b0010001111;
    cells[147] = 10'b0010001011;
    cells[148] = 10'b0010000111;
    cells[149] = 10'b0010000011;
    cells[150] = 10'b0001111111;
    cells[151] = 10'b0001111100;
    cells[152] = 10'b0001111000;
    cells[153] = 10'b0001110100;
    cells[154] = 10'b0001110000;
    cells[155] = 10'b0001101100;
    cells[156] = 10'b0001101000;
    cells[157] = 10'b0001100100;
    cells[158] = 10'b0001011111;
    cells[159] = 10'b0001011011;
    cells[160] = 10'b0001010111;
    cells[161] = 10'b0001010011;
    cells[162] = 10'b0001001111;
    cells[163] = 10'b0001001010;
    cells[164] = 10'b0001000110;
    cells[165] = 10'b0001000010;
    cells[166] = 10'b0000111101;
    cells[167] = 10'b0000111001;
    cells[168] = 10'b0000110101;
    cells[169] = 10'b0000110000;
    cells[170] = 10'b0000101100;
    cells[171] = 10'b0000101000;
    cells[172] = 10'b0000100011;
    cells[173] = 10'b0000011111;
    cells[174] = 10'b0000011010;
    cells[175] = 10'b0000010110;
    cells[176] = 10'b0000010001;
    cells[177] = 10'b0000001101;
    cells[178] = 10'b0000001000;
    cells[179] = 10'b0000000100;
    cells[180] = 10'b0000000000;
    cells[181] = 10'b1111111100;
    cells[182] = 10'b1111111000;
    cells[183] = 10'b1111110011;
    cells[184] = 10'b1111101111;
    cells[185] = 10'b1111101010;
    cells[186] = 10'b1111100110;
    cells[187] = 10'b1111100001;
    cells[188] = 10'b1111011101;
    cells[189] = 10'b1111011000;
    cells[190] = 10'b1111010100;
    cells[191] = 10'b1111010000;
    cells[192] = 10'b1111001011;
    cells[193] = 10'b1111000111;
    cells[194] = 10'b1111000011;
    cells[195] = 10'b1110111110;
    cells[196] = 10'b1110111010;
    cells[197] = 10'b1110110110;
    cells[198] = 10'b1110110001;
    cells[199] = 10'b1110101101;
    cells[200] = 10'b1110101001;
    cells[201] = 10'b1110100101;
    cells[202] = 10'b1110100001;
    cells[203] = 10'b1110011100;
    cells[204] = 10'b1110011000;
    cells[205] = 10'b1110010100;
    cells[206] = 10'b1110010000;
    cells[207] = 10'b1110001100;
    cells[208] = 10'b1110001000;
    cells[209] = 10'b1110000100;
    cells[210] = 10'b1110000000;
    cells[211] = 10'b1101111101;
    cells[212] = 10'b1101111001;
    cells[213] = 10'b1101110101;
    cells[214] = 10'b1101110001;
    cells[215] = 10'b1101101110;
    cells[216] = 10'b1101101010;
    cells[217] = 10'b1101100110;
    cells[218] = 10'b1101100011;
    cells[219] = 10'b1101011111;
    cells[220] = 10'b1101011100;
    cells[221] = 10'b1101011001;
    cells[222] = 10'b1101010101;
    cells[223] = 10'b1101010010;
    cells[224] = 10'b1101001111;
    cells[225] = 10'b1101001011;
    cells[226] = 10'b1101001000;
    cells[227] = 10'b1101000101;
    cells[228] = 10'b1101000010;
    cells[229] = 10'b1100111111;
    cells[230] = 10'b1100111100;
    cells[231] = 10'b1100111010;
    cells[232] = 10'b1100110111;
    cells[233] = 10'b1100110100;
    cells[234] = 10'b1100110001;
    cells[235] = 10'b1100101111;
    cells[236] = 10'b1100101100;
    cells[237] = 10'b1100101010;
    cells[238] = 10'b1100100111;
    cells[239] = 10'b1100100101;
    cells[240] = 10'b1100100011;
    cells[241] = 10'b1100100001;
    cells[242] = 10'b1100011110;
    cells[243] = 10'b1100011100;
    cells[244] = 10'b1100011010;
    cells[245] = 10'b1100011000;
    cells[246] = 10'b1100010111;
    cells[247] = 10'b1100010101;
    cells[248] = 10'b1100010011;
    cells[249] = 10'b1100010010;
    cells[250] = 10'b1100010000;
    cells[251] = 10'b1100001110;
    cells[252] = 10'b1100001101;
    cells[253] = 10'b1100001100;
    cells[254] = 10'b1100001010;
    cells[255] = 10'b1100001001;
    cells[256] = 10'b1100001000;
    cells[257] = 10'b1100000111;
    cells[258] = 10'b1100000110;
    cells[259] = 10'b1100000101;
    cells[260] = 10'b1100000100;
    cells[261] = 10'b1100000100;
    cells[262] = 10'b1100000011;
    cells[263] = 10'b1100000010;
    cells[264] = 10'b1100000010;
    cells[265] = 10'b1100000001;
    cells[266] = 10'b1100000001;
    cells[267] = 10'b1100000001;
    cells[268] = 10'b1100000001;
    cells[269] = 10'b1100000001;
    cells[270] = 10'b1100000000;
    cells[271] = 10'b1100000001;
    cells[272] = 10'b1100000001;
    cells[273] = 10'b1100000001;
    cells[274] = 10'b1100000001;
    cells[275] = 10'b1100000001;
    cells[276] = 10'b1100000010;
    cells[277] = 10'b1100000010;
    cells[278] = 10'b1100000011;
    cells[279] = 10'b1100000100;
    cells[280] = 10'b1100000100;
    cells[281] = 10'b1100000101;
    cells[282] = 10'b1100000110;
    cells[283] = 10'b1100000111;
    cells[284] = 10'b1100001000;
    cells[285] = 10'b1100001001;
    cells[286] = 10'b1100001010;
    cells[287] = 10'b1100001100;
    cells[288] = 10'b1100001101;
    cells[289] = 10'b1100001110;
    cells[290] = 10'b1100010000;
    cells[291] = 10'b1100010010;
    cells[292] = 10'b1100010011;
    cells[293] = 10'b1100010101;
    cells[294] = 10'b1100010111;
    cells[295] = 10'b1100011000;
    cells[296] = 10'b1100011010;
    cells[297] = 10'b1100011100;
    cells[298] = 10'b1100011110;
    cells[299] = 10'b1100100001;
    cells[300] = 10'b1100100011;
    cells[301] = 10'b1100100101;
    cells[302] = 10'b1100100111;
    cells[303] = 10'b1100101010;
    cells[304] = 10'b1100101100;
    cells[305] = 10'b1100101111;
    cells[306] = 10'b1100110001;
    cells[307] = 10'b1100110100;
    cells[308] = 10'b1100110111;
    cells[309] = 10'b1100111010;
    cells[310] = 10'b1100111100;
    cells[311] = 10'b1100111111;
    cells[312] = 10'b1101000010;
    cells[313] = 10'b1101000101;
    cells[314] = 10'b1101001000;
    cells[315] = 10'b1101001011;
    cells[316] = 10'b1101001111;
    cells[317] = 10'b1101010010;
    cells[318] = 10'b1101010101;
    cells[319] = 10'b1101011001;
    cells[320] = 10'b1101011100;
    cells[321] = 10'b1101011111;
    cells[322] = 10'b1101100011;
    cells[323] = 10'b1101100110;
    cells[324] = 10'b1101101010;
    cells[325] = 10'b1101101110;
    cells[326] = 10'b1101110001;
    cells[327] = 10'b1101110101;
    cells[328] = 10'b1101111001;
    cells[329] = 10'b1101111101;
    cells[330] = 10'b1110000001;
    cells[331] = 10'b1110000100;
    cells[332] = 10'b1110001000;
    cells[333] = 10'b1110001100;
    cells[334] = 10'b1110010000;
    cells[335] = 10'b1110010100;
    cells[336] = 10'b1110011000;
    cells[337] = 10'b1110011100;
    cells[338] = 10'b1110100001;
    cells[339] = 10'b1110100101;
    cells[340] = 10'b1110101001;
    cells[341] = 10'b1110101101;
    cells[342] = 10'b1110110001;
    cells[343] = 10'b1110110110;
    cells[344] = 10'b1110111010;
    cells[345] = 10'b1110111110;
    cells[346] = 10'b1111000011;
    cells[347] = 10'b1111000111;
    cells[348] = 10'b1111001011;
    cells[349] = 10'b1111010000;
    cells[350] = 10'b1111010100;
    cells[351] = 10'b1111011000;
    cells[352] = 10'b1111011101;
    cells[353] = 10'b1111100001;
    cells[354] = 10'b1111100110;
    cells[355] = 10'b1111101010;
    cells[356] = 10'b1111101111;
    cells[357] = 10'b1111110011;
    cells[358] = 10'b1111111000;
    cells[359] = 10'b1111111100;
    cells[360] = 0;
    cells[361] = 0;
    cells[362] = 0;
    cells[363] = 0;
    cells[364] = 0;
    cells[365] = 0;
    cells[366] = 0;
    cells[367] = 0;
    cells[368] = 0;
    cells[369] = 0;
    cells[370] = 0;
    cells[371] = 0;
    cells[372] = 0;
    cells[373] = 0;
    cells[374] = 0;
    cells[375] = 0;
    cells[376] = 0;
    cells[377] = 0;
    cells[378] = 0;
    cells[379] = 0;
    cells[380] = 0;
    cells[381] = 0;
    cells[382] = 0;
    cells[383] = 0;
    cells[384] = 0;
    cells[385] = 0;
    cells[386] = 0;
    cells[387] = 0;
    cells[388] = 0;
    cells[389] = 0;
    cells[390] = 0;
    cells[391] = 0;
    cells[392] = 0;
    cells[393] = 0;
    cells[394] = 0;
    cells[395] = 0;
    cells[396] = 0;
    cells[397] = 0;
    cells[398] = 0;
    cells[399] = 0;
    cells[400] = 0;
    cells[401] = 0;
    cells[402] = 0;
    cells[403] = 0;
    cells[404] = 0;
    cells[405] = 0;
    cells[406] = 0;
    cells[407] = 0;
    cells[408] = 0;
    cells[409] = 0;
    cells[410] = 0;
    cells[411] = 0;
    cells[412] = 0;
    cells[413] = 0;
    cells[414] = 0;
    cells[415] = 0;
    cells[416] = 0;
    cells[417] = 0;
    cells[418] = 0;
    cells[419] = 0;
    cells[420] = 0;
    cells[421] = 0;
    cells[422] = 0;
    cells[423] = 0;
    cells[424] = 0;
    cells[425] = 0;
    cells[426] = 0;
    cells[427] = 0;
    cells[428] = 0;
    cells[429] = 0;
    cells[430] = 0;
    cells[431] = 0;
    cells[432] = 0;
    cells[433] = 0;
    cells[434] = 0;
    cells[435] = 0;
    cells[436] = 0;
    cells[437] = 0;
    cells[438] = 0;
    cells[439] = 0;
    cells[440] = 0;
    cells[441] = 0;
    cells[442] = 0;
    cells[443] = 0;
    cells[444] = 0;
    cells[445] = 0;
    cells[446] = 0;
    cells[447] = 0;
    cells[448] = 0;
    cells[449] = 0;
    cells[450] = 0;
    cells[451] = 0;
    cells[452] = 0;
    cells[453] = 0;
    cells[454] = 0;
    cells[455] = 0;
    cells[456] = 0;
    cells[457] = 0;
    cells[458] = 0;
    cells[459] = 0;
    cells[460] = 0;
    cells[461] = 0;
    cells[462] = 0;
    cells[463] = 0;
    cells[464] = 0;
    cells[465] = 0;
    cells[466] = 0;
    cells[467] = 0;
    cells[468] = 0;
    cells[469] = 0;
    cells[470] = 0;
    cells[471] = 0;
    cells[472] = 0;
    cells[473] = 0;
    cells[474] = 0;
    cells[475] = 0;
    cells[476] = 0;
    cells[477] = 0;
    cells[478] = 0;
    cells[479] = 0;
    cells[480] = 0;
    cells[481] = 0;
    cells[482] = 0;
    cells[483] = 0;
    cells[484] = 0;
    cells[485] = 0;
    cells[486] = 0;
    cells[487] = 0;
    cells[488] = 0;
    cells[489] = 0;
    cells[490] = 0;
    cells[491] = 0;
    cells[492] = 0;
    cells[493] = 0;
    cells[494] = 0;
    cells[495] = 0;
    cells[496] = 0;
    cells[497] = 0;
    cells[498] = 0;
    cells[499] = 0;
    cells[500] = 0;
    cells[501] = 0;
    cells[502] = 0;
    cells[503] = 0;
    cells[504] = 0;
    cells[505] = 0;
    cells[506] = 0;
    cells[507] = 0;
    cells[508] = 0;
    cells[509] = 0;
    cells[510] = 0;
    cells[511] = 0;
end
endmodule

/*Produced by sfl2vl, IP ARCH, Inc. Sun Jul 14 18:45:28 2019
 Licensed to :EVALUATION USER*/
